LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY vga IS
PORT(
	CLOCK_50 :IN STD_LOGIC;
	VGA_HS:OUT STD_LOGIC;
	VGA_VS:OUT STD_LOGIC;
	VGA_BLANK:OUT STD_LOGIC;
	VGA_SYNC:OUT STD_LOGIC;
	VGA_CLK:OUT STD_LOGIC;
	VGA_R:OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	VGA_G:OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	VGA_B:OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END vga;

ARCHITECTURE main OF vga IS

COMPONENT vga_control IS
PORT(
	clk_50mz :IN STD_LOGIC;
	hsync:OUT STD_LOGIC;
	vsync:OUT STD_LOGIC;
	blank:OUT STD_LOGIC;
	sync:OUT STD_LOGIC;
	point_clk:OUT STD_LOGIC;
	x:OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
	y:OUT STD_LOGIC_VECTOR(10 DOWNTO 0)
	);
END COMPONENT;

COMPONENT graph_control IS
PORT(
	in_x: IN STD_LOGIC_VECTOR(10 DOWNTO 0);
	in_y: IN STD_LOGIC_VECTOR(10 DOWNTO 0);
	R:OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	G:OUT STD_LOGIC_VECTOR(9 DOWNTO 0);
	B:OUT STD_LOGIC_VECTOR(9 DOWNTO 0)
	);
END COMPONENT;

SIGNAL x: STD_LOGIC_VECTOR(10 DOWNTO 0);
SIGNAL y: STD_LOGIC_VECTOR(10 DOWNTO 0);

BEGIN

U1:vga_control PORT map(CLOCK_50, VGA_HS, VGA_VS, VGA_BLANK, VGA_SYNC, VGA_CLK, x, y);
U2:graph_control PORT map(x, y, VGA_R, VGA_G, VGA_B);

END main;
